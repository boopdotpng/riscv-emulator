module top #(
  parameter int Hello = 34
) (
  input logic [3:0] pause
);



endmodule
